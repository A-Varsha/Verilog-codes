`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 28.07.2025 07:56:23
// Design Name: 
// Module Name: summa_15
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module summa_15(
  input wire i0, i1, i2, i3,
  input wire S0, S1,
  output wire Y
);

  assign Y = S1 ? (S0 ? i3 : i2) : (S0 ? i1 : i0);

endmodule
